module OR_FOUR (a0,a1,a2,a3,y);
input logic a0,a1,a2,a3;
output logic y;
assign y = a0 | a1 | a2 | a3;
endmodule

